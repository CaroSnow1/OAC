library ieee;
use ieee.std_logic_1164.all;


entity registro is 
Port( clk : in std_logic;
		reset :  in std_logic;
		data_in: in std_logic_vector(2 downto 0); --LIGA
		data_out: out std_logic_vector(2 downto 0) --Edo
);
end registro;

architecture behavioral of registro is
	signal internal_value: std_logic_vector(2 downto 0):= B"000"; --Preguntar al profe
	begin
		process(clk, reset, data_in)
			begin 
			if reset = '0' then
				internal_value <= B"000";
			elsif rising_edge(clk) then 
				internal_value <= data_in;
			end if;
		end process;
		
	process(internal_value)
		begin
		data_out <= internal_value;
	end process;
end behavioral;
			